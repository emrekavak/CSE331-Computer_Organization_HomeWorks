module _32bitRight_shifter(res, inp1, inp0);
input [31:0]inp1;
input [31:0]inp0;
output[31:0]res;

wire [31:0]res00;
wire [31:0]res11;
wire [31:0]res22;
wire [31:0]res333;

_2x1mux _1(res00[0],inp1[1],inp1[0],inp0[0]);
_2x1mux _2(res00[1],inp1[2],inp1[1],inp0[0]);
_2x1mux _3(res00[2],inp1[3],inp1[2],inp0[0]);
_2x1mux _4(res00[3],inp1[4],inp1[3],inp0[0]);
_2x1mux _5(res00[4],inp1[5],inp1[4],inp0[0]);
_2x1mux _6(res00[5],inp1[6],inp1[5],inp0[0]);
_2x1mux _7(res00[6],inp1[7],inp1[6],inp0[0]);
_2x1mux _8(res00[7],inp1[8],inp1[7],inp0[0]);
_2x1mux _9(res00[8],inp1[9],inp1[8],inp0[0]);
_2x1mux _10(res00[9],inp1[10],inp1[9],inp0[0]);
_2x1mux _11(res00[10],inp1[11],inp1[10],inp0[0]);
_2x1mux _12(res00[11],inp1[12],inp1[11],inp0[0]);
_2x1mux _13(res00[12],inp1[13],inp1[12],inp0[0]);
_2x1mux _14(res00[13],inp1[14],inp1[13],inp0[0]);
_2x1mux _15(res00[14],inp1[15],inp1[14],inp0[0]);
_2x1mux _16(res00[15],inp1[16],inp1[15],inp0[0]);
_2x1mux _17(res00[16],inp1[17],inp1[16],inp0[0]);
_2x1mux _18(res00[17],inp1[18],inp1[17],inp0[0]);
_2x1mux _19(res00[18],inp1[19],inp1[18],inp0[0]);
_2x1mux _20(res00[19],inp1[20],inp1[19],inp0[0]);
_2x1mux _21(res00[20],inp1[21],inp1[20],inp0[0]);
_2x1mux _22(res00[21],inp1[22],inp1[21],inp0[0]);
_2x1mux _23(res00[22],inp1[23],inp1[22],inp0[0]);
_2x1mux _24(res00[23],inp1[24],inp1[23],inp0[0]);
_2x1mux _25(res00[24],inp1[25],inp1[24],inp0[0]);
_2x1mux _26(res00[25],inp1[26],inp1[25],inp0[0]);
_2x1mux _27(res00[26],inp1[27],inp1[26],inp0[0]);
_2x1mux _28(res00[27],inp1[28],inp1[27],inp0[0]);
_2x1mux _29(res00[28],inp1[29],inp1[28],inp0[0]);
_2x1mux _30(res00[29],inp1[30],inp1[29],inp0[0]);
_2x1mux _31(res00[30],inp1[31],inp1[30],inp0[0]);
_2x1mux _32(res00[31],inp1[31],inp1[31],inp0[0]);

_2x1mux _33(res11[0],res00[2],res00[0],inp0[1]);
_2x1mux _34(res11[1],res00[3],res00[1],inp0[1]);
_2x1mux _35(res11[2],res00[4],res00[2],inp0[1]);
_2x1mux _36(res11[3],res00[5],res00[3],inp0[1]);
_2x1mux _37(res11[4],res00[6],res00[4],inp0[1]);
_2x1mux _38(res11[5],res00[7],res00[5],inp0[1]);
_2x1mux _39(res11[6],res00[8],res00[6],inp0[1]);
_2x1mux _40(res11[7],res00[9],res00[7],inp0[1]);
_2x1mux _41(res11[8],res00[10],res00[8],inp0[1]);
_2x1mux _42(res11[9],res00[11],res00[9],inp0[1]);
_2x1mux _43(res11[10],res00[12],res00[10],inp0[1]);
_2x1mux _44(res11[11],res00[13],res00[11],inp0[1]);
_2x1mux _45(res11[12],res00[14],res00[12],inp0[1]);
_2x1mux _46(res11[13],res00[15],res00[13],inp0[1]);
_2x1mux _47(res11[14],res00[16],res00[14],inp0[1]);
_2x1mux _48(res11[15],res00[17],res00[15],inp0[1]);
_2x1mux _49(res11[16],res00[18],res00[16],inp0[1]);
_2x1mux _50(res11[17],res00[19],res00[17],inp0[1]);
_2x1mux _51(res11[18],res00[20],res00[18],inp0[1]);
_2x1mux _52(res11[19],res00[21],res00[19],inp0[1]);
_2x1mux _53(res11[20],res00[22],res00[20],inp0[1]);
_2x1mux _54(res11[21],res00[23],res00[21],inp0[1]);
_2x1mux _55(res11[22],res00[24],res00[22],inp0[1]);
_2x1mux _56(res11[23],res00[25],res00[23],inp0[1]);
_2x1mux _57(res11[24],res00[26],res00[24],inp0[1]);
_2x1mux _58(res11[25],res00[27],res00[25],inp0[1]);
_2x1mux _59(res11[26],res00[28],res00[26],inp0[1]);
_2x1mux _60(res11[27],res00[29],res00[27],inp0[1]);
_2x1mux _61(res11[28],res00[30],res00[28],inp0[1]);
_2x1mux _62(res11[29],res00[31],res00[29],inp0[1]);
_2x1mux _63(res11[30],res00[31],res00[30],inp0[1]);
_2x1mux _64(res11[31],res00[31],res00[31],inp0[1]);

_2x1mux _65(res22[0],res11[4],res11[0],inp0[2]);
_2x1mux _66(res22[1],res11[5],res11[1],inp0[2]);
_2x1mux _67(res22[2],res11[6],res11[2],inp0[2]);
_2x1mux _68(res22[3],res11[7],res11[3],inp0[2]);
_2x1mux _69(res22[4],res11[8],res11[4],inp0[2]);
_2x1mux _70(res22[5],res11[9],res11[5],inp0[2]);
_2x1mux _71(res22[6],res11[10],res11[6],inp0[2]);
_2x1mux _72(res22[7],res11[11],res11[7],inp0[2]);
_2x1mux _73(res22[8],res11[12],res11[8],inp0[2]);
_2x1mux _74(res22[9],res11[13],res11[9],inp0[2]);
_2x1mux _75(res22[10],res11[14],res11[10],inp0[2]);
_2x1mux _76(res22[11],res11[15],res11[11],inp0[2]);
_2x1mux _77(res22[12],res11[16],res11[12],inp0[2]);
_2x1mux _78(res22[13],res11[17],res11[13],inp0[2]);
_2x1mux _79(res22[14],res11[18],res11[14],inp0[2]);
_2x1mux _80(res22[15],res11[19],res11[15],inp0[2]);
_2x1mux _81(res22[16],res11[20],res11[16],inp0[2]);
_2x1mux _82(res22[17],res11[21],res11[17],inp0[2]);
_2x1mux _83(res22[18],res11[22],res11[18],inp0[2]);
_2x1mux _84(res22[19],res11[23],res11[19],inp0[2]);
_2x1mux _85(res22[20],res11[24],res11[20],inp0[2]);
_2x1mux _86(res22[21],res11[25],res11[21],inp0[2]);
_2x1mux _87(res22[22],res11[26],res11[22],inp0[2]);
_2x1mux _88(res22[23],res11[27],res11[23],inp0[2]);
_2x1mux _89(res22[24],res11[28],res11[24],inp0[2]);
_2x1mux _90(res22[25],res11[29],res11[25],inp0[2]);
_2x1mux _91(res22[26],res11[30],res11[26],inp0[2]);
_2x1mux _92(res22[27],res11[31],res11[27],inp0[2]);
_2x1mux _93(res22[28],res11[31],res11[28],inp0[2]);
_2x1mux _94(res22[29],res11[31],res11[29],inp0[2]);
_2x1mux _95(res22[30],res11[31],res11[30],inp0[2]);
_2x1mux _96(res22[31],res11[31],res11[31],inp0[2]);

_2x1mux _97(res333[0],res22[8],res22[0],inp0[3]);
_2x1mux _98(res333[1],res22[9],res22[1],inp0[3]);
_2x1mux _99(res333[2],res22[10],res22[2],inp0[3]);
_2x1mux _100(res333[3],res22[11],res22[3],inp0[3]);
_2x1mux _101(res333[4],res22[12],res22[4],inp0[3]);
_2x1mux _102(res333[5],res22[13],res22[5],inp0[3]);
_2x1mux _103(res333[6],res22[14],res22[6],inp0[3]);
_2x1mux _104(res333[7],res22[15],res22[7],inp0[3]);
_2x1mux _105(res333[8],res22[16],res22[8],inp0[3]);
_2x1mux _106(res333[9],res22[17],res22[9],inp0[3]);
_2x1mux _107(res333[10],res22[18],res22[10],inp0[3]);
_2x1mux _108(res333[11],res22[19],res22[11],inp0[3]);
_2x1mux _109(res333[12],res22[20],res22[12],inp0[3]);
_2x1mux _110(res333[13],res22[21],res22[13],inp0[3]);
_2x1mux _111(res333[14],res22[22],res22[14],inp0[3]);
_2x1mux _112(res333[15],res22[23],res22[15],inp0[3]);
_2x1mux _113(res333[16],res22[24],res22[16],inp0[3]);
_2x1mux _114(res333[17],res22[25],res22[17],inp0[3]);
_2x1mux _115(res333[18],res22[26],res22[18],inp0[3]);
_2x1mux _116(res333[19],res22[27],res22[19],inp0[3]);
_2x1mux _117(res333[20],res22[28],res22[20],inp0[3]);
_2x1mux _118(res333[21],res22[29],res22[21],inp0[3]);
_2x1mux _119(res333[22],res22[30],res22[22],inp0[3]);
_2x1mux _120(res333[23],res22[31],res22[23],inp0[3]);
_2x1mux _121(res333[24],res22[31],res22[24],inp0[3]);
_2x1mux _122(res333[25],res22[31],res22[25],inp0[3]);
_2x1mux _123(res333[26],res22[31],res22[26],inp0[3]);
_2x1mux _124(res333[27],res22[31],res22[27],inp0[3]);
_2x1mux _125(res333[28],res22[31],res22[28],inp0[3]);
_2x1mux _126(res333[29],res22[31],res22[29],inp0[3]);
_2x1mux _127(res333[30],res22[31],res22[30],inp0[3]);
_2x1mux _128(res333[31],res22[31],res22[31],inp0[3]);

_2x1mux _129(res[0],res333[16],res333[0],inp0[4]);
_2x1mux _130(res[1],res333[17],res333[1],inp0[4]);
_2x1mux _131(res[2],res333[18],res333[2],inp0[4]);
_2x1mux _132(res[3],res333[19],res333[3],inp0[4]);
_2x1mux _133(res[4],res333[20],res333[4],inp0[4]);
_2x1mux _134(res[5],res333[21],res333[5],inp0[4]);
_2x1mux _135(res[6],res333[22],res333[6],inp0[4]);
_2x1mux _136(res[7],res333[23],res333[7],inp0[4]);
_2x1mux _137(res[8],res333[24],res333[8],inp0[4]);
_2x1mux _138(res[9],res333[25],res333[9],inp0[4]);
_2x1mux _139(res[10],res333[26],res333[10],inp0[4]);
_2x1mux _140(res[11],res333[27],res333[11],inp0[4]);
_2x1mux _141(res[12],res333[28],res333[12],inp0[4]);
_2x1mux _142(res[13],res333[29],res333[13],inp0[4]);
_2x1mux _143(res[14],res333[30],res333[14],inp0[4]);
_2x1mux _144(res[15],res333[31],res333[15],inp0[4]);
_2x1mux _145(res[16],res333[31],res333[16],inp0[4]);
_2x1mux _146(res[17],res333[31],res333[17],inp0[4]);
_2x1mux _147(res[18],res333[31],res333[18],inp0[4]);
_2x1mux _148(res[19],res333[31],res333[19],inp0[4]);
_2x1mux _149(res[20],res333[31],res333[20],inp0[4]);
_2x1mux _150(res[21],res333[31],res333[21],inp0[4]);
_2x1mux _151(res[22],res333[31],res333[22],inp0[4]);
_2x1mux _152(res[23],res333[31],res333[23],inp0[4]);
_2x1mux _153(res[24],res333[31],res333[24],inp0[4]);
_2x1mux _154(res[25],res333[31],res333[25],inp0[4]);
_2x1mux _155(res[26],res333[31],res333[26],inp0[4]);
_2x1mux _156(res[27],res333[31],res333[27],inp0[4]);
_2x1mux _157(res[28],res333[31],res333[28],inp0[4]);
_2x1mux _158(res[29],res333[31],res333[29],inp0[4]);
_2x1mux _159(res[30],res333[31],res333[30],inp0[4]);
_2x1mux _160(res[31],res333[31],res333[31],inp0[4]);


endmodule