`define DELAY 10

module alu32_testbench();

reg [31:0] A;
reg [31:0] B;
reg[3:0] S;
wire [31:0] result;

alu32 test(result,A,B,S);

initial begin

A = 32'b11111111111111111111111111111111; 
B = 32'b11111111111111111111111111111111;
S= 3'b000;
#`DELAY;
A = 32'b10101010101010101010101010101010; 
B = 32'b01010101010101010101010101010101;
S= 3'b000;
#`DELAY;
A = 32'b10100010010000011111111111111111; 
B = 32'b10100010010000011111111111111111;
S= 3'b000;
#`DELAY;

//or
A = 32'b11111111111111111111111111111111; 
B = 32'b00000000000000000000000000000000;
S= 3'b001;
#`DELAY;
A = 32'b10101010101010101010101010101010; 
B = 32'b01010101010101010101010101010101;
S= 3'b001;
#`DELAY;
A = 32'b00111110111100011100011101011100; 
B = 32'b11000001000001100011100010100011;
S= 3'b001;
#`DELAY;

// adder
A = 32'b11111111111111111111111111111000; 
B = 32'b00000000000000000000000000000110;
S= 3'b010;
#`DELAY;
A = 32'b10000000000000000000000000000000; 
B = 32'b01000000000000001000000000000001;
S= 3'b010;
#`DELAY;
A = 32'b01010101010101010101010101010101; 
B = 32'b01010101010101010101010101010101;
S= 3'b010;
#`DELAY;

//xor
A = 32'b10101010101010101010101010101010; 
B = 32'b01010101010101010101010101010101;
S= 3'b011;
#`DELAY;
A = 32'b10101010101010101010101010101010; 
B = 32'b00000000000000000000000000000000;
S= 3'b011;
#`DELAY;
A = 32'b11111111111111111111111111111111; 
B = 32'b00000000000000000000000000000000;
S= 3'b011;
#`DELAY;

// subtrac
A = 32'b10101010101010101010101010101010; 
B = 32'b10101010101010101010101010101010;
S= 3'b100;
#`DELAY;
A = 32'b00000000000000000000000010000000; 
B = 32'b00000000000000000000000001010101;
S= 3'b100;
#`DELAY;
A = 32'b01111111111111111111111111111111; 
B = 32'b01010101010101010101010101010101;
S= 3'b100;
#`DELAY;

//right shift
A = 32'b10000000000000000000000000000000; 
B = 32'b00000000000000000000000000000011;
S= 3'b101;
#`DELAY;
A = 32'b10000000000000001111000000000000; 
B = 32'b00000000000000000000000000001100;
S= 3'b101;
#`DELAY;
A = 32'b10001110000000000000000000000000; 
B = 32'b00000000000000000000000000011111;
S= 3'b101;
#`DELAY;

//left shift
A = 32'b00000000000000000000000000000001; 
B = 32'b00000000000000000000000000111111;
S= 3'b110;
#`DELAY;
A = 32'b00000000000000000000000000011111; 
B = 32'b00000000000000000000000000000101;
S= 3'b110;
#`DELAY;
A = 32'b00000000000000000011111110000000; 
B = 32'b00000000000000000000000000001100;
S= 3'b110;
#`DELAY;

//nor
A = 32'b11111111111110001111111111111111; 
B = 32'b00000000000000000000000000000000;
S= 3'b111;
#`DELAY;
A = 32'b10101010101010101010101010101010; 
B = 32'b01010101010101010101010101010101;
S= 3'b111;
#`DELAY;
A = 32'b11001100110011001101100110011000; 
B = 32'b00000000000000000000000000000000;
S= 3'b111;
#`DELAY;

end


initial
begin
$monitor("A =%32b B=%32b \n S= %3b result-->%32b \n", A, B, S, result);
end
 
endmodule