module andop(andout,A,B);

input [31:0] A;
input [31:0] B;
output [31:0]andout;

and and0(andout[0],A[0],B[0]);
and and1(andout[1],A[1],B[1]);
and and2(andout[2],A[2],B[2]);
and and3(andout[3],A[3],B[3]);
and and4(andout[4],A[4],B[4]);
and and5(andout[5],A[5],B[5]);
and and6(andout[6],A[6],B[6]);
and and7(andout[7],A[7],B[7]);
and and8(andout[8],A[8],B[8]);
and and9(andout[9],A[9],B[9]);
and and10(andout[10],A[10],B[10]);
and and11(andout[11],A[11],B[11]);
and and12(andout[12],A[12],B[12]);
and and13(andout[13],A[13],B[13]);
and and14(andout[14],A[14],B[14]);
and and15(andout[15],A[15],B[15]);
and and16(andout[16],A[16],B[16]);
and and17(andout[17],A[17],B[17]);
and and18(andout[18],A[18],B[18]);
and and19(andout[19],A[19],B[19]);
and and20(andout[20],A[20],B[20]);
and and21(andout[21],A[21],B[21]);
and and22(andout[22],A[22],B[22]);
and and23(andout[23],A[23],B[23]);
and and24(andout[24],A[24],B[24]);
and and25(andout[25],A[25],B[25]);
and and26(andout[26],A[26],B[26]);
and and27(andout[27],A[27],B[27]);
and and28(andout[28],A[28],B[28]);
and and29(andout[29],A[29],B[29]);
and and30(andout[30],A[30],B[30]);
and and31(andout[31],A[31],B[31]);

endmodule