module _32bitLeft_shifter(reshifter, a1, b1);
input [31:0]a1;
input [31:0]b1;
output[31:0]reshifter;
wire [31:0]res0;
wire [31:0]res1;
wire [31:0]res2;
wire [31:0]res3;

_2x1mux _1(res0[0],1'b0,a1[0],b1[0]);
_2x1mux _2(res0[1],a1[0],a1[1],b1[0]);
_2x1mux _3(res0[2],a1[1],a1[2],b1[0]);
_2x1mux _4(res0[3],a1[2],a1[3],b1[0]);
_2x1mux _5(res0[4],a1[3],a1[4],b1[0]);
_2x1mux _6(res0[5],a1[4],a1[5],b1[0]);
_2x1mux _7(res0[6],a1[5],a1[6],b1[0]);
_2x1mux _8(res0[7],a1[6],a1[7],b1[0]);
_2x1mux _9(res0[8],a1[7],a1[8],b1[0]);
_2x1mux _10(res0[9],a1[8],a1[9],b1[0]);
_2x1mux _11(res0[10],a1[9],a1[10],b1[0]);
_2x1mux _12(res0[11],a1[10],a1[11],b1[0]);
_2x1mux _13(res0[12],a1[11],a1[12],b1[0]);
_2x1mux _14(res0[13],a1[12],a1[13],b1[0]);
_2x1mux _15(res0[14],a1[13],a1[14],b1[0]);
_2x1mux _16(res0[15],a1[14],a1[15],b1[0]);
_2x1mux _17(res0[16],a1[15],a1[16],b1[0]);
_2x1mux _18(res0[17],a1[16],a1[17],b1[0]);
_2x1mux _19(res0[18],a1[17],a1[18],b1[0]);
_2x1mux _20(res0[19],a1[18],a1[19],b1[0]);
_2x1mux _21(res0[20],a1[19],a1[20],b1[0]);
_2x1mux _22(res0[21],a1[20],a1[21],b1[0]);
_2x1mux _23(res0[22],a1[21],a1[22],b1[0]);
_2x1mux _24(res0[23],a1[22],a1[23],b1[0]);
_2x1mux _25(res0[24],a1[23],a1[24],b1[0]);
_2x1mux _26(res0[25],a1[24],a1[25],b1[0]);
_2x1mux _27(res0[26],a1[25],a1[26],b1[0]);
_2x1mux _28(res0[27],a1[26],a1[27],b1[0]);
_2x1mux _29(res0[28],a1[27],a1[28],b1[0]);
_2x1mux _30(res0[29],a1[28],a1[29],b1[0]);
_2x1mux _31(res0[30],a1[29],a1[30],b1[0]);
_2x1mux _32(res0[31],a1[30],a1[31],b1[0]);

_2x1mux _33(res1[0],1'b0,res0[0],b1[1]);
_2x1mux _34(res1[1],1'b0,res0[1],b1[1]);
_2x1mux _35(res1[2],res0[0],res0[2],b1[1]);
_2x1mux _36(res1[3],res0[1],res0[3],b1[1]);
_2x1mux _37(res1[4],res0[2],res0[4],b1[1]);
_2x1mux _38(res1[5],res0[3],res0[5],b1[1]);
_2x1mux _39(res1[6],res0[4],res0[6],b1[1]);
_2x1mux _40(res1[7],res0[5],res0[7],b1[1]);
_2x1mux _41(res1[8],res0[6],res0[8],b1[1]);
_2x1mux _42(res1[9],res0[7],res0[9],b1[1]);
_2x1mux _43(res1[10],res0[8],res0[10],b1[1]);
_2x1mux _44(res1[11],res0[9],res0[11],b1[1]);
_2x1mux _45(res1[12],res0[10],res0[12],b1[1]);
_2x1mux _46(res1[13],res0[11],res0[13],b1[1]);
_2x1mux _47(res1[14],res0[12],res0[14],b1[1]);
_2x1mux _48(res1[15],res0[13],res0[15],b1[1]);
_2x1mux _49(res1[16],res0[14],res0[16],b1[1]);
_2x1mux _50(res1[17],res0[15],res0[17],b1[1]);
_2x1mux _51(res1[18],res0[16],res0[18],b1[1]);
_2x1mux _52(res1[19],res0[17],res0[19],b1[1]);
_2x1mux _53(res1[20],res0[18],res0[20],b1[1]);
_2x1mux _54(res1[21],res0[19],res0[21],b1[1]);
_2x1mux _55(res1[22],res0[20],res0[22],b1[1]);
_2x1mux _56(res1[23],res0[21],res0[23],b1[1]);
_2x1mux _57(res1[24],res0[22],res0[24],b1[1]);
_2x1mux _58(res1[25],res0[23],res0[25],b1[1]);
_2x1mux _59(res1[26],res0[24],res0[26],b1[1]);
_2x1mux _60(res1[27],res0[25],res0[27],b1[1]);
_2x1mux _61(res1[28],res0[26],res0[28],b1[1]);
_2x1mux _62(res1[29],res0[27],res0[29],b1[1]);
_2x1mux _63(res1[30],res0[28],res0[30],b1[1]);
_2x1mux _64(res1[31],res0[29],res0[31],b1[1]);

_2x1mux _65(res2[0],1'b0,res1[0],b1[2]);
_2x1mux _66(res2[1],1'b0,res1[1],b1[2]);
_2x1mux _67(res2[2],1'b0,res1[2],b1[2]);
_2x1mux _68(res2[3],1'b0,res1[3],b1[2]);
_2x1mux _69(res2[4],res1[0],res1[4],b1[2]);
_2x1mux _70(res2[5],res1[1],res1[5],b1[2]);
_2x1mux _71(res2[6],res1[2],res1[6],b1[2]);
_2x1mux _72(res2[7],res1[3],res1[7],b1[2]);
_2x1mux _73(res2[8],res1[4],res1[8],b1[2]);
_2x1mux _74(res2[9],res1[5],res1[9],b1[2]);
_2x1mux _75(res2[10],res1[6],res1[10],b1[2]);
_2x1mux _76(res2[11],res1[7],res1[11],b1[2]);
_2x1mux _77(res2[12],res1[8],res1[12],b1[2]);
_2x1mux _78(res2[13],res1[9],res1[13],b1[2]);
_2x1mux _79(res2[14],res1[10],res1[14],b1[2]);
_2x1mux _80(res2[15],res1[11],res1[15],b1[2]);
_2x1mux _81(res2[16],res1[12],res1[16],b1[2]);
_2x1mux _82(res2[17],res1[13],res1[17],b1[2]);
_2x1mux _83(res2[18],res1[14],res1[18],b1[2]);
_2x1mux _84(res2[19],res1[15],res1[19],b1[2]);
_2x1mux _85(res2[20],res1[16],res1[20],b1[2]);
_2x1mux _86(res2[21],res1[17],res1[21],b1[2]);
_2x1mux _87(res2[22],res1[18],res1[22],b1[2]);
_2x1mux _88(res2[23],res1[19],res1[23],b1[2]);
_2x1mux _89(res2[24],res1[20],res1[24],b1[2]);
_2x1mux _90(res2[25],res1[21],res1[25],b1[2]);
_2x1mux _91(res2[26],res1[22],res1[26],b1[2]);
_2x1mux _92(res2[27],res1[23],res1[27],b1[2]);
_2x1mux _93(res2[28],res1[24],res1[28],b1[2]);
_2x1mux _94(res2[29],res1[25],res1[29],b1[2]);
_2x1mux _95(res2[30],res1[26],res1[30],b1[2]);
_2x1mux _96(res2[31],res1[27],res1[31],b1[2]);

_2x1mux _97(res3[0],1'b0,res2[0],b1[3]);
_2x1mux _98(res3[1],1'b0,res2[1],b1[3]);
_2x1mux _99(res3[2],1'b0,res2[2],b1[3]);
_2x1mux _100(res3[3],1'b0,res2[3],b1[3]);
_2x1mux _101(res3[4],1'b0,res2[4],b1[3]);
_2x1mux _102(res3[5],1'b0,res2[5],b1[3]);
_2x1mux _103(res3[6],1'b0,res2[6],b1[3]);
_2x1mux _104(res3[7],1'b0,res2[7],b1[3]);
_2x1mux _105(res3[8],res2[0],res2[8],b1[3]);
_2x1mux _106(res3[9],res2[1],res2[9],b1[3]);
_2x1mux _107(res3[10],res2[2],res2[10],b1[3]);
_2x1mux _108(res3[11],res2[3],res2[11],b1[3]);
_2x1mux _109(res3[12],res2[4],res2[12],b1[3]);
_2x1mux _110(res3[13],res2[5],res2[13],b1[3]);
_2x1mux _111(res3[14],res2[6],res2[14],b1[3]);
_2x1mux _112(res3[15],res2[7],res2[15],b1[3]);
_2x1mux _113(res3[16],res2[8],res2[16],b1[3]);
_2x1mux _114(res3[17],res2[9],res2[17],b1[3]);
_2x1mux _115(res3[18],res2[10],res2[18],b1[3]);
_2x1mux _116(res3[19],res2[11],res2[19],b1[3]);
_2x1mux _117(res3[20],res2[12],res2[20],b1[3]);
_2x1mux _118(res3[21],res2[13],res2[21],b1[3]);
_2x1mux _119(res3[22],res2[14],res2[22],b1[3]);
_2x1mux _120(res3[23],res2[15],res2[23],b1[3]);
_2x1mux _121(res3[24],res2[16],res2[24],b1[3]);
_2x1mux _122(res3[25],res2[17],res2[25],b1[3]);
_2x1mux _123(res3[26],res2[18],res2[26],b1[3]);
_2x1mux _124(res3[27],res2[19],res2[27],b1[3]);
_2x1mux _125(res3[28],res2[20],res2[28],b1[3]);
_2x1mux _126(res3[29],res2[21],res2[29],b1[3]);
_2x1mux _127(res3[30],res2[22],res2[30],b1[3]);
_2x1mux _128(res3[31],res2[23],res2[31],b1[3]);

_2x1mux _129(reshifter[0],1'b0,res3[0],b1[4]);
_2x1mux _130(reshifter[1],1'b0,res3[1],b1[4]);
_2x1mux _131(reshifter[2],1'b0,res3[2],b1[4]);
_2x1mux _132(reshifter[3],1'b0,res3[3],b1[4]);
_2x1mux _133(reshifter[4],1'b0,res3[4],b1[4]);
_2x1mux _134(reshifter[5],1'b0,res3[5],b1[4]);
_2x1mux _135(reshifter[6],1'b0,res3[6],b1[4]);
_2x1mux _136(reshifter[7],1'b0,res3[7],b1[4]);
_2x1mux _137(reshifter[8],1'b0,res3[8],b1[4]);
_2x1mux _138(reshifter[9],1'b0,res3[9],b1[4]);
_2x1mux _139(reshifter[10],1'b0,res3[10],b1[4]);
_2x1mux _140(reshifter[11],1'b0,res3[11],b1[4]);
_2x1mux _141(reshifter[12],1'b0,res3[12],b1[4]);
_2x1mux _142(reshifter[13],1'b0,res3[13],b1[4]);
_2x1mux _143(reshifter[14],1'b0,res3[14],b1[4]);
_2x1mux _144(reshifter[15],1'b0,res3[15],b1[4]);
_2x1mux _145(reshifter[16],res3[0],res3[16],b1[4]);
_2x1mux _146(reshifter[17],res3[1],res3[17],b1[4]);
_2x1mux _147(reshifter[18],res3[2],res3[18],b1[4]);
_2x1mux _148(reshifter[19],res3[3],res3[19],b1[4]);
_2x1mux _149(reshifter[20],res3[4],res3[20],b1[4]);
_2x1mux _150(reshifter[21],res3[5],res3[21],b1[4]);
_2x1mux _151(reshifter[22],res3[6],res3[22],b1[4]);
_2x1mux _152(reshifter[23],res3[7],res3[23],b1[4]);
_2x1mux _153(reshifter[24],res3[8],res3[24],b1[4]);
_2x1mux _154(reshifter[25],res3[9],res3[25],b1[4]);
_2x1mux _155(reshifter[26],res3[10],res3[26],b1[4]);
_2x1mux _156(reshifter[27],res3[11],res3[27],b1[4]);
_2x1mux _157(reshifter[28],res3[12],res3[28],b1[4]);
_2x1mux _158(reshifter[29],res3[13],res3[29],b1[4]);
_2x1mux _159(reshifter[30],res3[14],res3[30],b1[4]);
_2x1mux _160(reshifter[31],res3[15],res3[31],b1[4]);


endmodule